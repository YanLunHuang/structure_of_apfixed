`timescale 1 ns / 1 ps

module AESL_deadlock_detector (
    input reset,
    input clock);

    wire [0:0] proc_dep_vld_vec_0;
    reg [0:0] proc_dep_vld_vec_0_reg;
    wire [0:0] in_chan_dep_vld_vec_0;
    wire [2:0] in_chan_dep_data_vec_0;
    wire [0:0] token_in_vec_0;
    wire [0:0] out_chan_dep_vld_vec_0;
    wire [2:0] out_chan_dep_data_0;
    wire [0:0] token_out_vec_0;
    wire dl_detect_out_0;
    wire dep_chan_vld_1_0;
    wire [2:0] dep_chan_data_1_0;
    wire token_1_0;
    wire [1:0] proc_dep_vld_vec_1;
    reg [1:0] proc_dep_vld_vec_1_reg;
    wire [1:0] in_chan_dep_vld_vec_1;
    wire [5:0] in_chan_dep_data_vec_1;
    wire [1:0] token_in_vec_1;
    wire [1:0] out_chan_dep_vld_vec_1;
    wire [2:0] out_chan_dep_data_1;
    wire [1:0] token_out_vec_1;
    wire dl_detect_out_1;
    wire dep_chan_vld_0_1;
    wire [2:0] dep_chan_data_0_1;
    wire token_0_1;
    wire dep_chan_vld_2_1;
    wire [2:0] dep_chan_data_2_1;
    wire token_2_1;
    wire [0:0] proc_dep_vld_vec_2;
    reg [0:0] proc_dep_vld_vec_2_reg;
    wire [0:0] in_chan_dep_vld_vec_2;
    wire [2:0] in_chan_dep_data_vec_2;
    wire [0:0] token_in_vec_2;
    wire [0:0] out_chan_dep_vld_vec_2;
    wire [2:0] out_chan_dep_data_2;
    wire [0:0] token_out_vec_2;
    wire dl_detect_out_2;
    wire dep_chan_vld_1_2;
    wire [2:0] dep_chan_data_1_2;
    wire token_1_2;
    wire [2:0] dl_in_vec;
    wire dl_detect_out;
    wire [2:0] origin;
    wire token_clear;

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myproject$Block_proc_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myproject$Block_proc_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myproject$Block_proc_U0$ap_idle <= AESL_inst_myproject.Block_proc_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myproject.Block_proc_U0
    AESL_deadlock_detect_unit #(3, 0, 1, 1) AESL_deadlock_detect_unit_0 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_0),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_0),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_0),
        .token_in_vec(token_in_vec_0),
        .dl_detect_in(dl_detect_out),
        .origin(origin[0]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_0),
        .out_chan_dep_data(out_chan_dep_data_0),
        .token_out_vec(token_out_vec_0),
        .dl_detect_out(dl_in_vec[0]));

    assign proc_dep_vld_vec_0[0] = dl_detect_out ? proc_dep_vld_vec_0_reg[0] : (((AESL_inst_myproject.Block_proc_U0_ap_ready_count[0]) & AESL_inst_myproject.Block_proc_U0.ap_idle & ~(AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0_ap_ready_count[0])));
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_0_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_0_reg <= proc_dep_vld_vec_0;
        end
    end
    assign in_chan_dep_vld_vec_0[0] = dep_chan_vld_1_0;
    assign in_chan_dep_data_vec_0[2 : 0] = dep_chan_data_1_0;
    assign token_in_vec_0[0] = token_1_0;
    assign dep_chan_vld_0_1 = out_chan_dep_vld_vec_0[0];
    assign dep_chan_data_0_1 = out_chan_dep_data_0;
    assign token_0_1 = token_out_vec_0[0];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myproject$zeropad2d_cl_array_array_ap_fixed_256u_config4_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myproject$zeropad2d_cl_array_array_ap_fixed_256u_config4_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myproject$zeropad2d_cl_array_array_ap_fixed_256u_config4_U0$ap_idle <= AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0
    AESL_deadlock_detect_unit #(3, 1, 2, 2) AESL_deadlock_detect_unit_1 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_1),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_1),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_1),
        .token_in_vec(token_in_vec_1),
        .dl_detect_in(dl_detect_out),
        .origin(origin[1]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_1),
        .out_chan_dep_data(out_chan_dep_data_1),
        .token_out_vec(token_out_vec_1),
        .dl_detect_out(dl_in_vec[1]));

    assign proc_dep_vld_vec_1[0] = dl_detect_out ? proc_dep_vld_vec_1_reg[0] : (~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_0_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_1_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_2_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_3_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_4_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_5_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_6_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_7_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_8_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_9_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_10_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_11_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_12_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_13_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_14_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_15_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_16_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_17_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_18_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_19_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_20_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_21_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_22_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_23_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_24_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_25_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_26_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_27_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_28_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_29_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_30_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_31_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_32_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_33_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_34_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_35_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_36_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_37_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_38_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_39_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_40_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_41_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_42_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_43_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_44_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_45_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_46_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_47_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_48_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_49_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_50_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_51_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_52_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_53_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_54_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_55_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_56_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_57_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_58_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_59_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_60_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_61_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_62_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_63_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_64_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_65_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_66_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_67_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_68_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_69_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_70_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_71_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_72_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_73_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_74_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_75_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_76_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_77_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_78_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_79_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_80_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_81_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_82_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_83_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_84_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_85_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_86_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_87_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_88_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_89_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_90_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_91_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_92_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_93_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_94_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_95_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_96_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_97_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_98_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_99_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_100_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_101_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_102_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_103_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_104_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_105_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_106_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_107_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_108_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_109_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_110_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_111_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_112_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_113_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_114_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_115_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_116_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_117_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_118_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_119_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_120_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_121_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_122_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_123_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_124_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_125_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_126_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_127_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_128_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_129_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_130_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_131_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_132_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_133_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_134_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_135_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_136_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_137_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_138_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_139_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_140_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_141_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_142_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_143_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_144_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_145_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_146_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_147_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_148_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_149_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_150_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_151_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_152_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_153_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_154_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_155_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_156_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_157_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_158_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_159_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_160_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_161_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_162_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_163_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_164_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_165_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_166_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_167_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_168_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_169_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_170_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_171_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_172_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_173_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_174_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_175_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_176_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_177_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_178_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_179_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_180_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_181_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_182_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_183_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_184_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_185_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_186_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_187_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_188_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_189_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_190_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_191_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_192_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_193_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_194_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_195_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_196_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_197_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_198_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_199_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_200_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_201_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_202_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_203_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_204_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_205_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_206_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_207_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_208_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_209_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_210_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_211_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_212_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_213_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_214_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_215_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_216_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_217_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_218_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_219_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_220_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_221_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_222_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_223_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_224_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_225_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_226_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_227_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_228_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_229_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_230_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_231_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_232_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_233_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_234_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_235_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_236_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_237_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_238_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_239_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_240_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_241_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_242_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_243_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_244_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_245_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_246_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_247_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_248_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_249_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_250_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_251_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_252_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_253_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_254_V_blk_n | ~AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.res_V_data_255_V_blk_n | (~AESL_inst_myproject.start_for_conv_2d_cl_array_array_ap_fixed_256u_config2_U0_U.if_full_n & AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.ap_done));
    assign proc_dep_vld_vec_1[1] = dl_detect_out ? proc_dep_vld_vec_1_reg[1] : (((AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0_ap_ready_count[0]) & AESL_inst_myproject.zeropad2d_cl_array_array_ap_fixed_256u_config4_U0.ap_idle & ~(AESL_inst_myproject.Block_proc_U0_ap_ready_count[0])));
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_1_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_1_reg <= proc_dep_vld_vec_1;
        end
    end
    assign in_chan_dep_vld_vec_1[0] = dep_chan_vld_0_1;
    assign in_chan_dep_data_vec_1[2 : 0] = dep_chan_data_0_1;
    assign token_in_vec_1[0] = token_0_1;
    assign in_chan_dep_vld_vec_1[1] = dep_chan_vld_2_1;
    assign in_chan_dep_data_vec_1[5 : 3] = dep_chan_data_2_1;
    assign token_in_vec_1[1] = token_2_1;
    assign dep_chan_vld_1_2 = out_chan_dep_vld_vec_1[0];
    assign dep_chan_data_1_2 = out_chan_dep_data_1;
    assign token_1_2 = token_out_vec_1[0];
    assign dep_chan_vld_1_0 = out_chan_dep_vld_vec_1[1];
    assign dep_chan_data_1_0 = out_chan_dep_data_1;
    assign token_1_0 = token_out_vec_1[1];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myproject$conv_2d_cl_array_array_ap_fixed_256u_config2_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myproject$conv_2d_cl_array_array_ap_fixed_256u_config2_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myproject$conv_2d_cl_array_array_ap_fixed_256u_config2_U0$ap_idle <= AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0
    AESL_deadlock_detect_unit #(3, 2, 1, 1) AESL_deadlock_detect_unit_2 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_2),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_2),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_2),
        .token_in_vec(token_in_vec_2),
        .dl_detect_in(dl_detect_out),
        .origin(origin[2]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_2),
        .out_chan_dep_data(out_chan_dep_data_2),
        .token_out_vec(token_out_vec_2),
        .dl_detect_out(dl_in_vec[2]));

    assign proc_dep_vld_vec_2[0] = dl_detect_out ? proc_dep_vld_vec_2_reg[0] : (~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_0_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_1_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_2_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_3_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_4_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_5_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_6_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_7_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_8_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_9_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_10_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_11_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_12_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_13_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_14_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_15_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_16_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_17_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_18_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_19_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_20_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_21_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_22_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_23_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_24_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_25_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_26_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_27_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_28_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_29_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_30_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_31_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_32_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_33_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_34_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_35_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_36_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_37_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_38_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_39_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_40_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_41_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_42_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_43_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_44_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_45_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_46_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_47_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_48_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_49_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_50_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_51_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_52_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_53_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_54_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_55_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_56_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_57_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_58_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_59_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_60_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_61_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_62_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_63_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_64_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_65_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_66_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_67_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_68_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_69_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_70_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_71_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_72_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_73_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_74_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_75_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_76_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_77_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_78_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_79_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_80_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_81_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_82_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_83_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_84_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_85_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_86_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_87_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_88_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_89_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_90_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_91_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_92_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_93_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_94_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_95_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_96_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_97_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_98_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_99_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_100_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_101_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_102_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_103_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_104_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_105_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_106_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_107_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_108_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_109_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_110_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_111_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_112_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_113_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_114_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_115_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_116_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_117_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_118_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_119_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_120_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_121_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_122_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_123_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_124_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_125_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_126_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_127_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_128_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_129_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_130_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_131_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_132_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_133_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_134_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_135_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_136_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_137_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_138_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_139_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_140_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_141_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_142_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_143_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_144_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_145_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_146_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_147_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_148_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_149_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_150_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_151_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_152_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_153_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_154_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_155_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_156_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_157_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_158_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_159_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_160_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_161_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_162_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_163_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_164_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_165_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_166_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_167_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_168_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_169_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_170_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_171_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_172_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_173_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_174_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_175_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_176_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_177_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_178_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_179_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_180_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_181_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_182_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_183_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_184_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_185_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_186_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_187_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_188_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_189_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_190_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_191_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_192_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_193_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_194_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_195_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_196_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_197_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_198_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_199_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_200_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_201_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_202_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_203_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_204_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_205_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_206_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_207_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_208_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_209_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_210_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_211_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_212_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_213_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_214_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_215_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_216_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_217_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_218_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_219_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_220_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_221_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_222_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_223_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_224_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_225_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_226_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_227_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_228_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_229_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_230_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_231_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_232_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_233_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_234_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_235_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_236_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_237_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_238_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_239_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_240_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_241_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_242_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_243_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_244_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_245_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_246_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_247_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_248_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_249_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_250_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_251_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_252_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_253_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_254_V_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.data_V_data_255_V_blk_n | (~AESL_inst_myproject.start_for_conv_2d_cl_array_array_ap_fixed_256u_config2_U0_U.if_empty_n & (AESL_inst_myproject.conv_2d_cl_array_array_ap_fixed_256u_config2_U0.ap_ready | AESL_inst_myproject$conv_2d_cl_array_array_ap_fixed_256u_config2_U0$ap_idle)));
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_2_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_2_reg <= proc_dep_vld_vec_2;
        end
    end
    assign in_chan_dep_vld_vec_2[0] = dep_chan_vld_1_2;
    assign in_chan_dep_data_vec_2[2 : 0] = dep_chan_data_1_2;
    assign token_in_vec_2[0] = token_1_2;
    assign dep_chan_vld_2_1 = out_chan_dep_vld_vec_2[0];
    assign dep_chan_data_2_1 = out_chan_dep_data_2;
    assign token_2_1 = token_out_vec_2[0];


    AESL_deadlock_report_unit #(3) AESL_deadlock_report_unit_inst (
        .reset(reset),
        .clock(clock),
        .dl_in_vec(dl_in_vec),
        .dl_detect_out(dl_detect_out),
        .origin(origin),
        .token_clear(token_clear));

endmodule
